module imem(input  logic [31:0] a, output logic [31:0] rd);
  reg [31:0] ROM[255:0];
  initial begin
ROM[0]='hE04F000F;
ROM[1]='hE04F700F;
ROM[2]='hE28770FF;
ROM[3]='hE28770FF;
ROM[4]='hE28770FF;
ROM[5]='hE28020FF;
ROM[6]='hE5802804;
ROM[7]='hE5802804;
ROM[8]='hE2806050;
ROM[9]='hE080A00F;
ROM[10]='hEA000006;
ROM[11]='hE2806041;
ROM[12]='hE080A00F;
ROM[13]='hEA000003;
ROM[14]='hE2806049;
ROM[15]='hE080A00F;
ROM[16]='hEA000000;
ROM[17]='hEAFFFFFE;
ROM[18]='hE2861000;
ROM[19]='hE2513041;
ROM[20]='h0A000031;
ROM[21]='hE2513042;
ROM[22]='h0A000031;
ROM[23]='hE2513043;
ROM[24]='h0A000031;
ROM[25]='hE2513044;
ROM[26]='h0A000031;
ROM[27]='hE2513045;
ROM[28]='h0A000031;
ROM[29]='hE2513046;
ROM[30]='h0A000031;
ROM[31]='hE2513047;
ROM[32]='h0A000031;
ROM[33]='hE2513048;
ROM[34]='h0A000031;
ROM[35]='hE2513049;
ROM[36]='h0A000031;
ROM[37]='hE251304A;
ROM[38]='h0A000031;
ROM[39]='hE251304B;
ROM[40]='h0A000031;
ROM[41]='hE251304C;
ROM[42]='h0A000031;
ROM[43]='hE251304D;
ROM[44]='h0A000031;
ROM[45]='hE251304E;
ROM[46]='h0A000031;
ROM[47]='hE251304F;
ROM[48]='h0A000031;
ROM[49]='hE2513050;
ROM[50]='h0A000031;
ROM[51]='hE2513051;
ROM[52]='h0A000031;
ROM[53]='hE2513052;
ROM[54]='h0A000031;
ROM[55]='hE2513053;
ROM[56]='h0A000031;
ROM[57]='hE2513054;
ROM[58]='h0A000031;
ROM[59]='hE2513055;
ROM[60]='h0A000031;
ROM[61]='hE2513056;
ROM[62]='h0A000031;
ROM[63]='hE2513057;
ROM[64]='h0A000031;
ROM[65]='hE2513058;
ROM[66]='h0A000031;
ROM[67]='hE2513059;
ROM[68]='h0A000031;
ROM[69]='hE251305A;
ROM[70]='h0A000031;
ROM[71]='hE28010C4;
ROM[72]='hEA000031;
ROM[73]='hE28010F8;
ROM[74]='hEA00002F;
ROM[75]='hE28010FA;
ROM[76]='hEA00002D;
ROM[77]='hE28010E8;
ROM[78]='hEA00002B;
ROM[79]='hE2801080;
ROM[80]='hEA000029;
ROM[81]='hE28010F2;
ROM[82]='hEA000027;
ROM[83]='hE28010EC;
ROM[84]='hEA000025;
ROM[85]='hE28010F0;
ROM[86]='hEA000023;
ROM[87]='hE28010C0;
ROM[88]='hEA000021;
ROM[89]='hE28010F7;
ROM[90]='hEA00001F;
ROM[91]='hE28010EA;
ROM[92]='hEA00001D;
ROM[93]='hE28010F4;
ROM[94]='hEA00001B;
ROM[95]='hE28010CF;
ROM[96]='hEA000019;
ROM[97]='hE28010C8;
ROM[98]='hEA000017;
ROM[99]='hE28010EF;
ROM[100]='hEA000015;
ROM[101]='hE28010F6;
ROM[102]='hEA000013;
ROM[103]='hE28010FD;
ROM[104]='hEA000011;
ROM[105]='hE28010E4;
ROM[106]='hEA00000F;
ROM[107]='hE28010E0;
ROM[108]='hEA00000D;
ROM[109]='hE280108F;
ROM[110]='hEA00000B;
ROM[111]='hE28010E2;
ROM[112]='hEA000009;
ROM[113]='hE28010F1;
ROM[114]='hEA000007;
ROM[115]='hE28010E6;
ROM[116]='hEA000005;
ROM[117]='hE28010F9;
ROM[118]='hEA000003;
ROM[119]='hE28010FB;
ROM[120]='hEA000001;
ROM[121]='hE28010FC;
ROM[122]='hEAFFFFFF;
ROM[123]='hE2113008;
ROM[124]='hE080800F;
ROM[125]='h0A00001F;
ROM[126]='hE2113008;
ROM[127]='hE080800F;
ROM[128]='h1A000027;
ROM[129]='hE2113040;
ROM[130]='h0A000015;
ROM[131]='hE2113004;
ROM[132]='hE080800F;
ROM[133]='h0A000017;
ROM[134]='hE2113004;
ROM[135]='hE080800F;
ROM[136]='h1A00001F;
ROM[137]='hE2113020;
ROM[138]='h0A00000D;
ROM[139]='hE2113002;
ROM[140]='hE080800F;
ROM[141]='h0A00000F;
ROM[142]='hE2113002;
ROM[143]='hE080800F;
ROM[144]='h1A000017;
ROM[145]='hE2113010;
ROM[146]='h0A000005;
ROM[147]='hE2113001;
ROM[148]='hE080800F;
ROM[149]='h0A000007;
ROM[150]='hE2113001;
ROM[151]='hE080800F;
ROM[152]='h1A00000F;
ROM[153]='hE080900F;
ROM[154]='hEA00001C;
ROM[155]='hE080900F;
ROM[156]='hEA00001A;
ROM[157]='hE28AF000;
ROM[158]='hE2802001;
ROM[159]='hE5802800;
ROM[160]='hE5802800;
ROM[161]='hE080900F;
ROM[162]='hEA000014;
ROM[163]='hE2802000;
ROM[164]='hE5802800;
ROM[165]='hE5802800;
ROM[166]='hE080900F;
ROM[167]='hEA00000F;
ROM[168]='hE288F000;
ROM[169]='hE2802001;
ROM[170]='hE5802800;
ROM[171]='hE5802800;
ROM[172]='hE080900F;
ROM[173]='hEA000009;
ROM[174]='hE080900F;
ROM[175]='hEA000007;
ROM[176]='hE080900F;
ROM[177]='hEA000005;
ROM[178]='hE2802000;
ROM[179]='hE5802800;
ROM[180]='hE5802800;
ROM[181]='hE080900F;
ROM[182]='hEA000000;
ROM[183]='hE288F000;
ROM[184]='hE04F400F;
ROM[185]='hE2445001;
ROM[186]='hE0555007;
ROM[187]='h7AFFFFFD;
ROM[188]='hE289F000;
  end
  assign rd = ROM[a[31:2]];
endmodule